module ula();
	
endmodule 